library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity instr_mem is
    port
    (
        clk: in std_logic;
        rd_addr: in std_logic_vector (31 downto 0);
        rd_data: out std_logic_vector (31 downto 0);
        wr_en: in std_logic;
        wr_addr: in std_logic_vector (31 downto 0);
        wr_data: in std_logic_vector (31 downto 0)
    );
end instr_mem;

architecture behav of instr_mem is
    type MEMORY is array (0 to 1023) of std_logic_vector (31 downto 0);

    signal mem : MEMORY := (
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000026",
        x"00000826",
        x"00001026",
        x"00001826",
        x"00002026",
        x"00002826",
        x"00003026",
        x"00003826",
        x"00004026",
        x"00004826",
        x"00005026",
        x"00005826",
        x"00006026",
        x"00006826",
        x"00007026",
        x"00007826",
        x"00008026",
        x"00008826",
        x"00009026",
        x"00009826",
        x"0000a026",
        x"0000a826",
        x"0000b026",
        x"0000b826",
        x"0000c026",
        x"0000c826",
        x"0000d026",
        x"0000d826",
        x"0000e026",
        x"0000e826",
        x"0000f026",
        x"0000f826",
        x"20150000",
        x"20170100",
        x"20160180",
        x"20100800",
        x"20141000",
        x"201d4000",
        x"20134000",
        x"20114010",
        x"20125000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"2001000b",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"ae610000",
        x"20080010",
        x"22090000",
        x"201a007f",
        x"201b0040",
        x"2001000c",
        x"a1200000",
        x"a1200001",
        x"a13a0002",
        x"a13b0003",
        x"a13a0004",
        x"a1200005",
        x"a1200006",
        x"a1210007",
        x"ad200008",
        x"2129000c",
        x"2108ffff",
        x"2101ffff",
        x"0020082a",
        x"1020ffef",
        x"00000000",
        x"00000000",
        x"00000000",
        x"2001000c",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"ae610000",
        x"20080040",
        x"22490000",
        x"2001ffff",
        x"ad200000",
        x"ad200004",
        x"ad200008",
        x"ad20000c",
        x"ad210010",
        x"ad210014",
        x"ad200018",
        x"ad20001c",
        x"21290020",
        x"2108ffff",
        x"2101ffff",
        x"0020082a",
        x"1020fff2",
        x"00000000",
        x"00000000",
        x"00000000",
        x"20010002",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"ae610000",
        x"8e280004",
        x"00000000",
        x"00000000",
        x"00000000",
        x"1100fffb",
        x"00000000",
        x"00000000",
        x"00000000",
        x"8e280000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00084902",
        x"3108000f",
        x"00000000",
        x"00000000",
        x"20010008",
        x"1121002b",
        x"00000000",
        x"00000000",
        x"00000000",
        x"20010009",
        x"11210070",
        x"00000000",
        x"00000000",
        x"00000000",
        x"2001000a",
        x"11210141",
        x"00000000",
        x"00000000",
        x"00000000",
        x"2001000b",
        x"1121015e",
        x"00000000",
        x"00000000",
        x"00000000",
        x"2001000c",
        x"1121020b",
        x"00000000",
        x"00000000",
        x"00000000",
        x"2001000d",
        x"11210224",
        x"00000000",
        x"00000000",
        x"00000000",
        x"2001000e",
        x"11210235",
        x"00000000",
        x"00000000",
        x"00000000",
        x"2001000f",
        x"112102a2",
        x"00000000",
        x"00000000",
        x"00000000",
        x"200400f1",
        x"100002df",
        x"00000000",
        x"00000000",
        x"00000000",
        x"20010003",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"ae610000",
        x"8e2a0004",
        x"00000000",
        x"00000000",
        x"00000000",
        x"1140fffb",
        x"00000000",
        x"00000000",
        x"00000000",
        x"8e2a0000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"8e210004",
        x"00000000",
        x"00000000",
        x"00000000",
        x"1020fffb",
        x"00000000",
        x"00000000",
        x"00000000",
        x"8e210000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"20090040",
        x"00125821",
        x"816c0001",
        x"00000000",
        x"00000000",
        x"00000000",
        x"018ad02a",
        x"014cd82a",
        x"035bd027",
        x"335a0001",
        x"13400015",
        x"00000000",
        x"00000000",
        x"00000000",
        x"816c0005",
        x"00000000",
        x"00000000",
        x"00000000",
        x"0188d02a",
        x"010cd82a",
        x"035bd027",
        x"335a0001",
        x"13400009",
        x"00000000",
        x"00000000",
        x"00000000",
        x"200c0010",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"a16c0000",
        x"216b0020",
        x"2129ffff",
        x"2121ffff",
        x"0020082a",
        x"1020ffdd",
        x"00000000",
        x"00000000",
        x"00000000",
        x"1000ff76",
        x"00000000",
        x"00000000",
        x"00000000",
        x"20010004",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"ae610000",
        x"8e2a0004",
        x"00000000",
        x"00000000",
        x"00000000",
        x"1140fffb",
        x"00000000",
        x"00000000",
        x"00000000",
        x"8e2a0000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"8e2d0004",
        x"00000000",
        x"00000000",
        x"00000000",
        x"11a0fffb",
        x"00000000",
        x"00000000",
        x"00000000",
        x"8e2d0000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"11a0ffb5",
        x"00000000",
        x"00000000",
        x"00000000",
        x"20090040",
        x"00125821",
        x"816c0000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"20010000",
        x"11810025",
        x"00000000",
        x"00000000",
        x"00000000",
        x"216b0020",
        x"2129ffff",
        x"2121ffff",
        x"0020082a",
        x"1020fff2",
        x"00000000",
        x"00000000",
        x"00000000",
        x"20090040",
        x"00125821",
        x"816c0000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"20010001",
        x"11810012",
        x"00000000",
        x"00000000",
        x"00000000",
        x"216b0020",
        x"2129ffff",
        x"2121ffff",
        x"0020082a",
        x"1020fff2",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00125821",
        x"200100aa",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"ae610000",
        x"200c0008",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"a16c0000",
        x"200c000c",
        x"71886002",
        x"01906020",
        x"00000000",
        x"00000000",
        x"00000000",
        x"818e0002",
        x"818f0004",
        x"81980003",
        x"00000000",
        x"00000000",
        x"00000000",
        x"71ae0802",
        x"702f0802",
        x"2002007f",
        x"00581022",
        x"00181820",
        x"70411002",
        x"00021502",
        x"02a2d020",
        x"83420000",
        x"70611802",
        x"00031d02",
        x"02a3d820",
        x"83630000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"a1620002",
        x"a1630003",
        x"a16a0001",
        x"a1680005",
        x"a16d0006",
        x"818e0000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"200d0018",
        x"71ae6802",
        x"01b46820",
        x"20010009",
        x"0101d02a",
        x"0028d82a",
        x"035bd027",
        x"335a0001",
        x"13400010",
        x"00000000",
        x"00000000",
        x"00000000",
        x"2001007f",
        x"11c1000b",
        x"00000000",
        x"00000000",
        x"00000000",
        x"200d0018",
        x"71aa6802",
        x"01b46820",
        x"21ad0c00",
        x"00000000",
        x"00000000",
        x"00000000",
        x"81aa0001",
        x"8dae0008",
        x"8daf000c",
        x"8db80010",
        x"8db90014",
        x"00000000",
        x"ad6e0010",
        x"ad6f0014",
        x"ad780018",
        x"ad79001c",
        x"8dae0004",
        x"81af0000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"ad6e000c",
        x"a16f0004",
        x"00000000",
        x"00000000",
        x"00000000",
        x"818d0007",
        x"8d8e0008",
        x"00000000",
        x"00000000",
        x"00000000",
        x"71ae0802",
        x"00010943",
        x"303a00ff",
        x"00010a03",
        x"0141d820",
        x"03771020",
        x"80430001",
        x"80420000",
        x"00000000",
        x"3044000f",
        x"00042080",
        x"00021102",
        x"3065000f",
        x"00052880",
        x"00031902",
        x"02c40820",
        x"8c240000",
        x"02c50820",
        x"8c250000",
        x"00000000",
        x"00000000",
        x"00442006",
        x"00652806",
        x"00a41022",
        x"000210c2",
        x"705a1002",
        x"00021142",
        x"00441020",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"ad620008",
        x"20080020",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"a1680000",
        x"1000fea0",
        x"00000000",
        x"00000000",
        x"00000000",
        x"20010005",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"ae610000",
        x"8e280004",
        x"00000000",
        x"00000000",
        x"00000000",
        x"1100fffb",
        x"00000000",
        x"00000000",
        x"00000000",
        x"8e280000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"8e280004",
        x"00000000",
        x"00000000",
        x"00000000",
        x"1100fffb",
        x"00000000",
        x"00000000",
        x"00000000",
        x"8e280000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"1000fe7e",
        x"00000000",
        x"00000000",
        x"00000000",
        x"20010006",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"ae610000",
        x"8e290004",
        x"00000000",
        x"00000000",
        x"00000000",
        x"1120fffb",
        x"00000000",
        x"00000000",
        x"00000000",
        x"8e290000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"8e2a0004",
        x"00000000",
        x"00000000",
        x"00000000",
        x"1140fffb",
        x"00000000",
        x"00000000",
        x"00000000",
        x"8e2a0000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"200b000c",
        x"71685802",
        x"01705820",
        x"20010006",
        x"11210016",
        x"00000000",
        x"00000000",
        x"00000000",
        x"20010007",
        x"11210032",
        x"00000000",
        x"00000000",
        x"00000000",
        x"2001000a",
        x"11210036",
        x"00000000",
        x"00000000",
        x"00000000",
        x"2001000b",
        x"1121003a",
        x"00000000",
        x"00000000",
        x"00000000",
        x"1000fe45",
        x"00000000",
        x"00000000",
        x"00000000",
        x"816c0005",
        x"00000000",
        x"00000000",
        x"00000000",
        x"0180d02a",
        x"000cd82a",
        x"035bd027",
        x"335a0001",
        x"1340fe39",
        x"00000000",
        x"00000000",
        x"00000000",
        x"816c0006",
        x"00000000",
        x"00000000",
        x"00000000",
        x"0180d02a",
        x"000cd82a",
        x"035bd027",
        x"335a0001",
        x"1340fe2d",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"a16a0007",
        x"1000fe24",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"a16a0002",
        x"10000015",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"a16a0003",
        x"1000000c",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"a16a0004",
        x"10000003",
        x"00000000",
        x"00000000",
        x"00000000",
        x"81690002",
        x"816a0003",
        x"816c0004",
        x"200e0040",
        x"224b0000",
        x"816d0005",
        x"00000000",
        x"00000000",
        x"00000000",
        x"01a8d02a",
        x"010dd82a",
        x"035bd027",
        x"335a0001",
        x"13400023",
        x"00000000",
        x"00000000",
        x"00000000",
        x"816d0000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"20010001",
        x"11a1001a",
        x"00000000",
        x"00000000",
        x"00000000",
        x"816d0006",
        x"00000000",
        x"00000000",
        x"00000000",
        x"71a90802",
        x"702c0802",
        x"2002007f",
        x"004a1022",
        x"000a1820",
        x"70411002",
        x"00021502",
        x"02a2d020",
        x"83420000",
        x"70611802",
        x"00031d02",
        x"02a3d820",
        x"83630000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"a1620002",
        x"a1630003",
        x"216b0020",
        x"21ceffff",
        x"21c1ffff",
        x"0020082a",
        x"1020ffcf",
        x"00000000",
        x"00000000",
        x"00000000",
        x"1000fdcc",
        x"00000000",
        x"00000000",
        x"00000000",
        x"20010007",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"ae610000",
        x"8e290004",
        x"00000000",
        x"00000000",
        x"00000000",
        x"1120fffb",
        x"00000000",
        x"00000000",
        x"00000000",
        x"8e290000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"200a000c",
        x"71485002",
        x"01505020",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"a1490000",
        x"1000fdae",
        x"00000000",
        x"00000000",
        x"00000000",
        x"20010008",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"ae610000",
        x"8e280004",
        x"00000000",
        x"00000000",
        x"00000000",
        x"1100fffb",
        x"00000000",
        x"00000000",
        x"00000000",
        x"8e280000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"1000fd98",
        x"00000000",
        x"00000000",
        x"00000000",
        x"20010009",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"ae610000",
        x"8e290004",
        x"00000000",
        x"00000000",
        x"00000000",
        x"1120fffb",
        x"00000000",
        x"00000000",
        x"00000000",
        x"8e290000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"8e2a0004",
        x"00000000",
        x"00000000",
        x"00000000",
        x"1140fffb",
        x"00000000",
        x"00000000",
        x"00000000",
        x"8e2a0000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"000a51c0",
        x"012a4825",
        x"2129e000",
        x"200b000c",
        x"71685802",
        x"01705820",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"ad690008",
        x"816e0007",
        x"200a0040",
        x"224c0000",
        x"818d0005",
        x"00000000",
        x"00000000",
        x"00000000",
        x"01a8d02a",
        x"010dd82a",
        x"035bd027",
        x"335a0001",
        x"13400031",
        x"00000000",
        x"00000000",
        x"00000000",
        x"818d0000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"20010001",
        x"11a10028",
        x"00000000",
        x"00000000",
        x"00000000",
        x"818d0001",
        x"00000000",
        x"00000000",
        x"00000000",
        x"712e0802",
        x"00010943",
        x"303a00ff",
        x"00010a03",
        x"01a1d820",
        x"03771020",
        x"80430001",
        x"80420000",
        x"00000000",
        x"3044000f",
        x"00042080",
        x"00021102",
        x"3065000f",
        x"00052880",
        x"00031902",
        x"02c40820",
        x"8c240000",
        x"02c50820",
        x"8c250000",
        x"00000000",
        x"00000000",
        x"00442006",
        x"00652806",
        x"00a41022",
        x"000210c2",
        x"705a1002",
        x"00021142",
        x"00441020",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"ad820008",
        x"218c0020",
        x"214affff",
        x"2141ffff",
        x"0020082a",
        x"1020ffc1",
        x"00000000",
        x"00000000",
        x"00000000",
        x"1000fd26",
        x"00000000",
        x"00000000",
        x"00000000",
        x"2001000a",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"ae610000",
        x"00144020",
        x"20091800",
        x"8e2a0004",
        x"00000000",
        x"00000000",
        x"00000000",
        x"1140fffb",
        x"00000000",
        x"00000000",
        x"00000000",
        x"8e2a0000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"a10a0000",
        x"00090982",
        x"34210080",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"a2610000",
        x"21080001",
        x"2129ffff",
        x"2121ffff",
        x"0020082a",
        x"1020ffe3",
        x"00000000",
        x"00000000",
        x"00000000",
        x"8e280004",
        x"00000000",
        x"00000000",
        x"00000000",
        x"1100fffb",
        x"00000000",
        x"00000000",
        x"00000000",
        x"8e280000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"200400f2",
        x"200100f7",
        x"0101d02a",
        x"0028d82a",
        x"035bd027",
        x"335a0001",
        x"13400007",
        x"00000000",
        x"00000000",
        x"00000000",
        x"1000fcaf",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"00000000",
        x"ae640000",
        x"1000ffff",
        x"00000000",
        x"00000000",
        x"00000000",
        others => (others => '0')
    );
begin
    process (clk)
    begin
        if (rising_edge(clk)) then
            rd_data <= mem(to_integer(unsigned(rd_addr(11 downto 2))));
            if (wr_en = '1') then
                mem(to_integer(unsigned(wr_addr(11 downto 2)))) <= wr_data;
            end if;
        end if;
    end process;
end architecture;
